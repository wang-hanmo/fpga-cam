module fpga_cam_tb;

endmodule